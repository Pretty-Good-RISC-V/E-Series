import PGRV::*;

import MachineInformation::*;
import MachineISA::*;
import MachineStatus::*;

export MachineInformation::*, MachineISA::*, MachineStatus::*;
